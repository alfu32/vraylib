@[translated]
module main
